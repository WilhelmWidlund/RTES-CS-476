
module soc_system (
	accelerator_0_conduit_end_readdata,
	clk_clk,
	reset_reset_n);	

	output	[7:0]	accelerator_0_conduit_end_readdata;
	input		clk_clk;
	input		reset_reset_n;
endmodule
