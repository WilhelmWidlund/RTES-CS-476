-- #############################################################################
-- DE1_SoC_top_level.vhd
--
-- BOARD         : DE1-SoC from Terasic
-- Author        : Sahand Kashani-Akhavan from Terasic documentation
-- Revision      : 1.4
-- Creation date : 04/02/2015
--
-- Syntax Rule : GROUP_NAME_N[bit]
--
-- GROUP  : specify a particular interface (ex: SDR_)
-- NAME   : signal name (ex: CONFIG, D, ...)
-- bit    : signal index
-- _N     : to specify an active-low signal
-- #############################################################################

library ieee;
use ieee.std_logic_1164.all;

entity DE1_SoC_top_level is
    port(
        -- ADC
--        ADC_CS_n         : out   std_logic;
--        ADC_DIN          : out   std_logic;
--        ADC_DOUT         : in    std_logic;
--        ADC_SCLK         : out   std_logic;

        -- Audio
        AUD_ADCDAT       : in    std_logic;
        AUD_ADCLRCK      : inout std_logic;
        AUD_BCLK         : inout std_logic;
        AUD_DACDAT       : out   std_logic;
        AUD_DACLRCK      : inout std_logic;
        AUD_XCK          : out   std_logic;

        -- CLOCK
        CLOCK_50         : in    std_logic;
--        CLOCK2_50        : in    std_logic;
--        CLOCK3_50        : in    std_logic;
--        CLOCK4_50        : in    std_logic;

        -- SDRAM
        DRAM_ADDR        : out   std_logic_vector(12 downto 0);
        DRAM_BA          : out   std_logic_vector(1 downto 0);
        DRAM_CAS_N       : out   std_logic;
        DRAM_CKE         : out   std_logic;
        DRAM_CLK         : out   std_logic;
        DRAM_CS_N        : out   std_logic;
        DRAM_DQ          : inout std_logic_vector(15 downto 0);
        DRAM_LDQM        : out   std_logic;
        DRAM_RAS_N       : out   std_logic;
        DRAM_UDQM        : out   std_logic;
        DRAM_WE_N        : out   std_logic;

        -- I2C for Audio and Video-In
        FPGA_I2C_SCLK    : out   std_logic;
        FPGA_I2C_SDAT    : inout std_logic;

        -- SEG7
        HEX0_N           : out   std_logic_vector(6 downto 0);
        HEX1_N           : out   std_logic_vector(6 downto 0);
        HEX2_N           : out   std_logic_vector(6 downto 0);
        HEX3_N           : out   std_logic_vector(6 downto 0);
        HEX4_N           : out   std_logic_vector(6 downto 0);
        HEX5_N           : out   std_logic_vector(6 downto 0);

        -- IR
--        IRDA_RXD         : in    std_logic;
--        IRDA_TXD         : out   std_logic;

        -- KEY_N
        KEY_N            : in    std_logic_vector(3 downto 0);

        -- LED
        LEDR             : out   std_logic_vector(9 downto 0);

        -- PS2
--        PS2_CLK          : inout std_logic;
--        PS2_CLK2         : inout std_logic;
--        PS2_DAT          : inout std_logic;
--        PS2_DAT2         : inout std_logic;

        -- SW
        SW               : in    std_logic_vector(9 downto 0)

        -- Video-In
--        TD_CLK27         : inout std_logic;
--        TD_DATA          : out   std_logic_vector(7 downto 0);
--        TD_HS            : out   std_logic;
--        TD_RESET_N       : out   std_logic;
--        TD_VS            : out   std_logic;

        -- VGA
--        VGA_B            : out   std_logic_vector(7 downto 0);
--        VGA_BLANK_N      : out   std_logic;
--        VGA_CLK          : out   std_logic;
--        VGA_G            : out   std_logic_vector(7 downto 0);
--        VGA_HS           : out   std_logic;
--        VGA_R            : out   std_logic_vector(7 downto 0);
--        VGA_SYNC_N       : out   std_logic;
--        VGA_VS           : out   std_logic;

        -- GPIO_0
--        GPIO_0           : inout std_logic_vector(35 downto 0);

        -- GPIO_1
--        GPIO_1           : inout std_logic_vector(35 downto 0);

        -- HPS
--        HPS_CONV_USB_N   : inout std_logic;
--        HPS_DDR3_ADDR    : out   std_logic_vector(14 downto 0);
--        HPS_DDR3_BA      : out   std_logic_vector(2 downto 0);
--        HPS_DDR3_CAS_N   : out   std_logic;
--        HPS_DDR3_CK_N    : out   std_logic;
--        HPS_DDR3_CK_P    : out   std_logic;
--        HPS_DDR3_CKE     : out   std_logic;
--        HPS_DDR3_CS_N    : out   std_logic;
--        HPS_DDR3_DM      : out   std_logic_vector(3 downto 0);
--        HPS_DDR3_DQ      : inout std_logic_vector(31 downto 0);
--        HPS_DDR3_DQS_N   : inout std_logic_vector(3 downto 0);
--        HPS_DDR3_DQS_P   : inout std_logic_vector(3 downto 0);
--        HPS_DDR3_ODT     : out   std_logic;
--        HPS_DDR3_RAS_N   : out   std_logic;
--        HPS_DDR3_RESET_N : out   std_logic;
--        HPS_DDR3_RZQ     : in    std_logic;
--        HPS_DDR3_WE_N    : out   std_logic;
--        HPS_ENET_GTX_CLK : out   std_logic;
--        HPS_ENET_INT_N   : inout std_logic;
--        HPS_ENET_MDC     : out   std_logic;
--        HPS_ENET_MDIO    : inout std_logic;
--        HPS_ENET_RX_CLK  : in    std_logic;
--        HPS_ENET_RX_DATA : in    std_logic_vector(3 downto 0);
--        HPS_ENET_RX_DV   : in    std_logic;
--        HPS_ENET_TX_DATA : out   std_logic_vector(3 downto 0);
--        HPS_ENET_TX_EN   : out   std_logic;
--        HPS_FLASH_DATA   : inout std_logic_vector(3 downto 0);
--        HPS_FLASH_DCLK   : out   std_logic;
--        HPS_FLASH_NCSO   : out   std_logic;
--        HPS_GSENSOR_INT  : inout std_logic;
--        HPS_I2C_CONTROL  : inout std_logic;
--        HPS_I2C1_SCLK    : inout std_logic;
--        HPS_I2C1_SDAT    : inout std_logic;
--        HPS_I2C2_SCLK    : inout std_logic;
--        HPS_I2C2_SDAT    : inout std_logic;
--        HPS_KEY_N        : inout std_logic;
--        HPS_LED          : inout std_logic;
--        HPS_LTC_GPIO     : inout std_logic;
--        HPS_SD_CLK       : out   std_logic;
--        HPS_SD_CMD       : inout std_logic;
--        HPS_SD_DATA      : inout std_logic_vector(3 downto 0);
--        HPS_SPIM_CLK     : out   std_logic;
--        HPS_SPIM_MISO    : in    std_logic;
--        HPS_SPIM_MOSI    : out   std_logic;
--        HPS_SPIM_SS      : inout std_logic;
--        HPS_UART_RX      : in    std_logic;
--        HPS_UART_TX      : out   std_logic;
--        HPS_USB_CLKOUT   : in    std_logic;
--        HPS_USB_DATA     : inout std_logic_vector(7 downto 0);
--        HPS_USB_DIR      : in    std_logic;
--        HPS_USB_NXT      : in    std_logic;
--        HPS_USB_STP      : out   std_logic
    );
end entity DE1_SoC_top_level;

architecture rtl of DE1_SoC_top_level is

component soc_system is
		port (
			clk_clk                                        : in    std_logic                     := 'X';             -- clk
			in_switches_export                             : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			out_led_export                                 : out   std_logic_vector(9 downto 0);                    -- export
			pll_shared_outclk2_clk                         : out   std_logic;                                        -- clk
			reset_reset_n                                  : in    std_logic                     := 'X';             -- reset_n
			sdram_controller_shared_wire_addr              : out   std_logic_vector(12 downto 0);                    -- addr
			sdram_controller_shared_wire_ba                : out   std_logic_vector(1 downto 0);                     -- ba
			sdram_controller_shared_wire_cas_n             : out   std_logic;                                        -- cas_n
			sdram_controller_shared_wire_cke               : out   std_logic;                                        -- cke
			sdram_controller_shared_wire_cs_n              : out   std_logic;                                        -- cs_n
			sdram_controller_shared_wire_dq                : inout std_logic_vector(31 downto 0) := (others => 'X'); -- dq
			sdram_controller_shared_wire_dqm               : out   std_logic_vector(3 downto 0);                     -- dqm
			sdram_controller_shared_wire_ras_n             : out   std_logic;                                        -- ras_n
			sdram_controller_shared_wire_we_n              : out   std_logic;                                        -- we_n
			sysaudio_audio_core_external_interface_ADCDAT  : in    std_logic                     := 'X';             -- ADCDAT
			sysaudio_audio_core_external_interface_ADCLRCK : in    std_logic                     := 'X';             -- ADCLRCK
			sysaudio_audio_core_external_interface_BCLK    : in    std_logic                     := 'X';             -- BCLK
			sysaudio_audio_core_external_interface_DACDAT  : out   std_logic;                                        -- DACDAT
			sysaudio_audio_core_external_interface_DACLRCK : in    std_logic                     := 'X';             -- DACLRCK
			sysaudio_av_config_external_interface_SDAT     : inout std_logic                     := 'X';             -- SDAT
			sysaudio_av_config_external_interface_SCLK     : out   std_logic;                                        -- SCLK
			pio_1st_7seg_external_connection_export        : out   std_logic_vector(13 downto 0);                    -- export
			pio_2nd_7seg_external_connection_export        : out   std_logic_vector(13 downto 0);                    -- export
			pio_3rd_7seg_external_connection_export        : out   std_logic_vector(13 downto 0)                     -- export
		);
	end component soc_system;

begin

u0 : component soc_system
		port map (
			clk_clk                                        => CLOCK_50,                                        --                                    clk.clk
			in_switches_export                             => SW(7 downto 0),                             --                            in_switches.export
			out_led_export                                 => LEDR(9 downto 0),                                 --                                out_led.export
			pll_shared_outclk2_clk                         => DRAM_CLK,                         --                     pll_shared_outclk2.clk
			reset_reset_n                                  => KEY_N(0),                                  --                                  reset.reset_n
			sdram_controller_shared_wire_addr              => DRAM_ADDR,              --           sdram_controller_shared_wire.addr
			sdram_controller_shared_wire_ba                => DRAM_BA,                --                                       .ba
			sdram_controller_shared_wire_cas_n             => DRAM_CAS_N,             --                                       .cas_n
			sdram_controller_shared_wire_cke               => DRAM_CKE,               --                                       .cke
			sdram_controller_shared_wire_cs_n              => DRAM_CS_N,              --                                       .cs_n
			sdram_controller_shared_wire_dq                => DRAM_DQ,                --                                       .dq
			sdram_controller_shared_wire_dqm(1)            => DRAM_UDQM,               --                                       .dqm(1)
			sdram_controller_shared_wire_dqm(0)            => DRAM_LDQM,               --                                       .dqm(0)
			sdram_controller_shared_wire_ras_n             => DRAM_RAS_N,             --                                       .ras_n
			sdram_controller_shared_wire_we_n              => DRAM_WE_N,              --                                       .we_n
			
			-- Audio
			-- TODO: Connected these just by name, seems straightforward enough
        --AUD_ADCDAT       : in    std_logic;
        --AUD_ADCLRCK      : inout std_logic;
        --AUD_BCLK         : inout std_logic;
        --AUD_DACDAT       : out   std_logic;
        --AUD_DACLRCK      : inout std_logic;
        -- TODO: This guy goes where??? Is it like that this guy is not used because of the whole Audio Clock IP thing???
		  --AUD_XCK          : out   std_logic;
			
			sysaudio_audio_core_external_interface_ADCDAT  => AUD_ADCDAT,  -- sysaudio_audio_core_external_interface.ADCDAT
			sysaudio_audio_core_external_interface_ADCLRCK => AUD_ADCLRCK, --                                       .ADCLRCK
			sysaudio_audio_core_external_interface_BCLK    => AUD_BCLK,    --                                       .BCLK
			sysaudio_audio_core_external_interface_DACDAT  => AUD_DACDAT,  --                                       .DACDAT
			sysaudio_audio_core_external_interface_DACLRCK => AUD_DACLRCK, --                                       .DACLRCK
			
			-- I2C for Audio and Video-In
			-- TODO: These seem to have similar names, so I made these connections. However I have no idea really...
        --FPGA_I2C_SCLK    : out   std_logic;
        --FPGA_I2C_SDAT    : inout std_logic;
			
			sysaudio_av_config_external_interface_SDAT     => FPGA_I2C_SDAT,     --  sysaudio_av_config_external_interface.SDAT
			sysaudio_av_config_external_interface_SCLK     => FPGA_I2C_SCLK,     --                                       .SCLK
			
			-- TODO: Which order does this correspond to??? 
			pio_1st_7seg_external_connection_export(13 downto 7)        => HEX0_N,        --       pio_1st_7seg_external_connection.export
			pio_1st_7seg_external_connection_export(6 downto 0)        => HEX1_N,
			pio_2nd_7seg_external_connection_export(13 downto 7)        => HEX2_N,        --       pio_2nd_7seg_external_connection.export
			pio_2nd_7seg_external_connection_export(6 downto 0)        => HEX3_N,
			pio_3rd_7seg_external_connection_export(13 downto 7)        => HEX4_N,        --       pio_3rd_7seg_external_connection.export
			pio_3rd_7seg_external_connection_export(6 downto 0)        => HEX5_N      
		);
		
		
end;
